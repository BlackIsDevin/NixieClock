////////////////////////////////////////////////////////////////////////////////
// File: Testbench-ClockStateStorage.v
// Author: BlackIsDevin (https://github.com/BlackIsDevin)
// Creation Date: 3/27/2021‏‎
// Target Devices: Mimas A7 Revision V3 Development Board 
//
// Description: This module is intended to test and verify the functionality of
// the ClockStateStorage module.
////////////////////////////////////////////////////////////////////////////////

module TestbenchClockStateStorage(

);

endmodule