////////////////////////////////////////////////////////////////////////////////
// File: NixieSignalGeneration.v
// Author: BlackIsDevin (https://github.com/BlackIsDevin)
// Creation Date: 3/23/2021‏‎
// Target Devices: Mimas A7 Revision V3 Development Board 
//
// Description: This module takes in the value of the clock state, and generates
// the appropriate signals to drive the nixie tubes.
////////////////////////////////////////////////////////////////////////////////