////////////////////////////////////////////////////////////////////////////////
// File: InputHandler.v
// Author: BlackIsDevin (https://github.com/BlackIsDevin)
// Creation Date: 3/23/2021‏‎
// Target Devices: Mimas A7 Revision V3 Development Board 
//
// Description: This module parses the user input (buttons and dip switches) 
// and generates signals for the ClockStateStorage module to interpret.
////////////////////////////////////////////////////////////////////////////////