////////////////////////////////////////////////////////////////////////////////
// File: NixieClockTopModule.v
// Author: BlackIsDevin (https://github.com/BlackIsDevin)
// Creation Date: 3/23/2021‏‎
// Target Devices: Mimas A7 Revision V3 Development Board 
//
// Description: This module links together all the underlying modules for the
// NixieClock project and exposes inputs and outputs for the FPGA and any
// testbench modules.
////////////////////////////////////////////////////////////////////////////////